module booth (X, Y, Z,en);
       input signed [15:0] X, Y;
   input en;
       output signed [31:0] Z;
       reg signed [31:0] Z;
       reg [1:0] temp;
       integer i;
       reg E1;
       reg [15:0] Y1;
       always @ (X, Y,en)
       begin
       Z = 32'd0;
       E1 = 1'd0;
       for (i = 0; i < 16; i = i + 1)
       begin
       temp = {X[i], E1};
      
           //The above statement is catenation
      
       Y1 = - Y;
      
           //Y1 is the 2� complement of Y
      
       case (temp)
       2'd2 : Z [31 : 15] = Z [31 : 15] + Y1;
       2'd1 : Z [31 : 15] = Z [31 : 15] + Y;
       default : begin end
       endcase
       Z = Z >> 1;
       /*The above statement is a logical shift of one position to
           the right*/
      
       Z[31] = Z[30];
       /*The above two statements perform arithmetic shift where
       the sign of the number is preserved after the shift. */
      
       E1 = X[i];
           end
       if (Y == 16'd32)
      
       /*If Y = 1000; then according to our code,
       Y1 = 1000 (-8 not 8, because Y1 is 4 bits only).
       The statement sum = - sum adjusts the answer.*/
      
           begin
               Z = - Z;
           end
      
       end
      
       endmodule
